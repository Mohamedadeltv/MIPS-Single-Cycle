`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:56:17 03/17/2021 
// Design Name: 
// Module Name:    thirdsection 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module thirdsection(
    input [31:0] A,
    input [31:0] B,
    input [3:0] OPERATION,
    output ZERO,
    output [31:0] C
    );


endmodule
